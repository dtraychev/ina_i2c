// module ina_top #(
//     parameters
// )(
//     port_list
// );
    
// endmodule
